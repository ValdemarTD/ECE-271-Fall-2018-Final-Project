module NES_Decoder(
  input logic Sig, clk, Latch,
  output logic [4:0]
);
